// Generator : SpinalHDL v1.3.8    git head : 57d97088b91271a094cebad32ed86479199955df
// Date      : 06/04/2021, 01:42:40
// Component : testMatrix


module testMatrix (
      input   clk,
      input   reset);
  wire [8:0] _zz_23_;
  wire [8:0] _zz_24_;
  wire [8:0] _zz_25_;
  wire [8:0] _zz_26_;
  wire [8:0] _zz_27_;
  wire [8:0] _zz_28_;
  wire [8:0] _zz_29_;
  wire [8:0] _zz_30_;
  wire [8:0] _zz_31_;
  wire [8:0] _zz_32_;
  wire [8:0] _zz_33_;
  wire [8:0] _zz_34_;
  reg [7:0] m1_mat_0_0;
  reg [7:0] m1_mat_0_1;
  reg [7:0] m1_mat_1_0;
  reg [7:0] m1_mat_1_1;
  reg [7:0] m2_mat_0_0;
  reg [7:0] m2_mat_0_1;
  reg [7:0] m2_mat_1_0;
  reg [7:0] m2_mat_1_1;
  reg [7:0] m3_mat_0_0;
  reg [7:0] m3_mat_0_1;
  reg [7:0] m3_mat_1_0;
  reg [7:0] m3_mat_1_1;
  reg [8:0] m4_mat_0_0;
  reg [8:0] m4_mat_0_1;
  reg [8:0] m4_mat_1_0;
  reg [8:0] m4_mat_1_1;
  reg [8:0] _zz_1_;
  reg [8:0] _zz_2_;
  reg [8:0] _zz_3_;
  reg [8:0] _zz_4_;
  reg [15:0] m1_mul_Matrix2D_0_0_0;
  wire [7:0] _zz_5_;
  reg [15:0] m1_mul_Matrix2D_0_0_1;
  wire [7:0] _zz_6_;
  reg [8:0] _zz_7_;
  reg [15:0] m1_mul_Matrix2D_0_1_0;
  wire [7:0] _zz_8_;
  reg [15:0] m1_mul_Matrix2D_0_1_1;
  wire [7:0] _zz_9_;
  reg [8:0] _zz_10_;
  reg [8:0] m5_mat_0_0;
  reg [8:0] m5_mat_0_1;
  reg [8:0] m5_mat_1_0;
  reg [8:0] m5_mat_1_1;
  reg [15:0] m1_mul_Matrix2D_0_0_0_1_;
  wire [7:0] _zz_11_;
  reg [15:0] m1_mul_Matrix2D_0_0_1_1_;
  wire [7:0] _zz_12_;
  reg [8:0] _zz_13_;
  reg [15:0] m1_mul_Matrix2D_0_1_0_1_;
  wire [7:0] _zz_14_;
  reg [15:0] m1_mul_Matrix2D_0_1_1_1_;
  wire [7:0] _zz_15_;
  reg [8:0] _zz_16_;
  reg [15:0] m1_mul_Matrix2D_1_0_0;
  wire [7:0] _zz_17_;
  reg [15:0] m1_mul_Matrix2D_1_0_1;
  wire [7:0] _zz_18_;
  reg [8:0] _zz_19_;
  reg [15:0] m1_mul_Matrix2D_1_1_0;
  wire [7:0] _zz_20_;
  reg [15:0] m1_mul_Matrix2D_1_1_1;
  wire [7:0] _zz_21_;
  reg [8:0] _zz_22_;
  assign _zz_23_ = {_zz_5_[7],_zz_5_};
  assign _zz_24_ = {_zz_6_[7],_zz_6_};
  assign _zz_25_ = {_zz_8_[7],_zz_8_};
  assign _zz_26_ = {_zz_9_[7],_zz_9_};
  assign _zz_27_ = {_zz_11_[7],_zz_11_};
  assign _zz_28_ = {_zz_12_[7],_zz_12_};
  assign _zz_29_ = {_zz_14_[7],_zz_14_};
  assign _zz_30_ = {_zz_15_[7],_zz_15_};
  assign _zz_31_ = {_zz_17_[7],_zz_17_};
  assign _zz_32_ = {_zz_18_[7],_zz_18_};
  assign _zz_33_ = {_zz_20_[7],_zz_20_};
  assign _zz_34_ = {_zz_21_[7],_zz_21_};
  assign _zz_5_ = m1_mul_Matrix2D_0_0_0[15 : 8];
  assign _zz_6_ = m1_mul_Matrix2D_0_0_1[15 : 8];
  assign _zz_8_ = m1_mul_Matrix2D_0_1_0[15 : 8];
  assign _zz_9_ = m1_mul_Matrix2D_0_1_1[15 : 8];
  assign _zz_11_ = m1_mul_Matrix2D_0_0_0_1_[15 : 8];
  assign _zz_12_ = m1_mul_Matrix2D_0_0_1_1_[15 : 8];
  assign _zz_14_ = m1_mul_Matrix2D_0_1_0_1_[15 : 8];
  assign _zz_15_ = m1_mul_Matrix2D_0_1_1_1_[15 : 8];
  assign _zz_17_ = m1_mul_Matrix2D_1_0_0[15 : 8];
  assign _zz_18_ = m1_mul_Matrix2D_1_0_1[15 : 8];
  assign _zz_20_ = m1_mul_Matrix2D_1_1_0[15 : 8];
  assign _zz_21_ = m1_mul_Matrix2D_1_1_1[15 : 8];
  always @ (posedge clk) begin
    m2_mat_0_0 <= m2_mat_0_1;
    m2_mat_1_0 <= m2_mat_1_1;
    m2_mat_0_1 <= m2_mat_0_0;
    m2_mat_1_1 <= m2_mat_1_0;
    m3_mat_0_0 <= m1_mat_0_0;
    m3_mat_0_1 <= m1_mat_0_1;
    m3_mat_1_0 <= m2_mat_1_0;
    m3_mat_1_1 <= m2_mat_1_1;
    m1_mat_0_0 <= m1_mat_1_0;
    m1_mat_0_1 <= m1_mat_1_1;
    m1_mat_1_0 <= m1_mat_0_0;
    m1_mat_1_1 <= m1_mat_0_1;
    m1_mul_Matrix2D_0_0_0 <= ($signed(m1_mat_0_0) * $signed(m2_mat_0_0));
    m1_mul_Matrix2D_0_0_1 <= ($signed(m1_mat_0_1) * $signed(m2_mat_1_0));
    _zz_7_ <= ($signed(_zz_23_) + $signed(_zz_24_));
    _zz_1_ <= _zz_7_;
    m1_mul_Matrix2D_0_1_0 <= ($signed(m1_mat_0_0) * $signed(m2_mat_0_1));
    m1_mul_Matrix2D_0_1_1 <= ($signed(m1_mat_0_1) * $signed(m2_mat_1_1));
    _zz_10_ <= ($signed(_zz_25_) + $signed(_zz_26_));
    _zz_2_ <= _zz_10_;
    _zz_3_ <= _zz_1_;
    _zz_4_ <= _zz_2_;
    m4_mat_0_0 <= _zz_1_;
    m4_mat_0_1 <= _zz_2_;
    m4_mat_1_0 <= _zz_3_;
    m4_mat_1_1 <= _zz_4_;
    m1_mul_Matrix2D_0_0_0_1_ <= ($signed(m1_mat_0_0) * $signed(m2_mat_0_0));
    m1_mul_Matrix2D_0_0_1_1_ <= ($signed(m1_mat_0_1) * $signed(m2_mat_1_0));
    _zz_13_ <= ($signed(_zz_27_) + $signed(_zz_28_));
    m5_mat_0_0 <= _zz_13_;
    m1_mul_Matrix2D_0_1_0_1_ <= ($signed(m1_mat_0_0) * $signed(m2_mat_0_1));
    m1_mul_Matrix2D_0_1_1_1_ <= ($signed(m1_mat_0_1) * $signed(m2_mat_1_1));
    _zz_16_ <= ($signed(_zz_29_) + $signed(_zz_30_));
    m5_mat_0_1 <= _zz_16_;
    m1_mul_Matrix2D_1_0_0 <= ($signed(m1_mat_1_0) * $signed(m2_mat_0_0));
    m1_mul_Matrix2D_1_0_1 <= ($signed(m1_mat_1_1) * $signed(m2_mat_1_0));
    _zz_19_ <= ($signed(_zz_31_) + $signed(_zz_32_));
    m5_mat_1_0 <= _zz_19_;
    m1_mul_Matrix2D_1_1_0 <= ($signed(m1_mat_1_0) * $signed(m2_mat_0_1));
    m1_mul_Matrix2D_1_1_1 <= ($signed(m1_mat_1_1) * $signed(m2_mat_1_1));
    _zz_22_ <= ($signed(_zz_33_) + $signed(_zz_34_));
    m5_mat_1_1 <= _zz_22_;
  end

endmodule

